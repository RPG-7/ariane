/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 860;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h0a0d2165_6e6f6420,
        64'h00000000_00206567,
        64'h616d6920_746f6f62,
        64'h20676e69_79706f63,
        64'h00000000_00000009,
        64'h3a656d61_6e090a0d,
        64'h00093a73_65747562,
        64'h69727474_61090a0d,
        64'h00000009_3a61626c,
        64'h20747361_6c090a0d,
        64'h0000093a_61626c20,
        64'h74737269_66090a0d,
        64'h00000000_00000000,
        64'h09202020_20203a64,
        64'h69756720_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_00000000,
        64'h093a6469_75672065,
        64'h70797420_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20747067,
        64'h00000009_20203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20657a69_73090a0d,
        64'h00000009_3a736569,
        64'h72746e65_206e6f69,
        64'h74697472_61702072,
        64'h65626d75_6e090a0d,
        64'h00000009_2020203a,
        64'h61626c20_73656972,
        64'h746e6520_6e6f6974,
        64'h69747261_70090a0d,
        64'h00093a61_646c2070,
        64'h756b6361_62090a0d,
        64'h00000000_00000000,
        64'h093a6162_6c20746e,
        64'h65727275_63090a0d,
        64'h00000009_3a646576,
        64'h72657365_72090a0d,
        64'h00093a72_65646165,
        64'h685f6372_63090a0d,
        64'h00000000_00000909,
        64'h3a657a69_73090a0d,
        64'h00000009_3a6e6f69,
        64'h73697665_72090a0d,
        64'h0000093a_65727574,
        64'h616e6769_73090a0d,
        64'h00000000_003a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20747067,
        64'h0000203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_63206473,
        64'h00000000_0000000a,
        64'h0d216465_6c696166,
        64'h20647261_63204453,
        64'h00000000_0000000a,
        64'h0d216465_7a696c61,
        64'h6974696e_69206473,
        64'h00000000_0a0d676e,
        64'h69746978_65202e2e,
        64'h2e647320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f63,
        64'h00000000_0000002e,
        64'h0000000a_0d202e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e69,
        64'h00000031_34646d63,
        64'h00000035_35646d63,
        64'h00000000_30646d63,
        64'h00000020_3a206573,
        64'h6e6f7073_65720920,
        64'h00000000_0020646e,
        64'h616d6d6f_63204453,
        64'h00000000_203f3f79,
        64'h74706d65_20746f6e,
        64'h206f6669_66207872,
        64'h00000000_00000a0d,
        64'h2164657a_696c6169,
        64'h74696e69_20495053,
        64'h00000000_00007830,
        64'h203a7375_74617473,
        64'h00000000_00000a0d,
        64'h49505320_74696e69,
        64'h00000a0d_21646c72,
        64'h6f57206f_6c6c6548,
        64'h00000000_00006564,
        64'h6f6d2d79_6870006f,
        64'h69646d2d_7361682c,
        64'h786e6c78_006c616e,
        64'h7265746e_692d6573,
        64'h752c786e_6c780067,
        64'h6e6f702d_676e6970,
        64'h2d78742c_786e6c78,
        64'h00687464_69772d64,
        64'h692d6978_612d732c,
        64'h786e6c78_00676e6f,
        64'h702d676e_69702d78,
        64'h722c786e_6c780065,
        64'h636e6174_736e692c,
        64'h786e6c78_006f6964,
        64'h6d2d6564_756c636e,
        64'h692c786e_6c78006b,
        64'h63616270_6f6f6c2d,
        64'h6c616e72_65746e69,
        64'h2d656475_6c636e69,
        64'h2c786e6c_78007372,
        64'h65666675_622d6c61,
        64'h626f6c67_2d656475,
        64'h6c636e69_2c786e6c,
        64'h78007865_6c707564,
        64'h2c786e6c_7800656c,
        64'h646e6168_2d796870,
        64'h00737365_72646461,
        64'h2d63616d_2d6c6163,
        64'h6f6c0070_772d656c,
        64'h62617369_64007365,
        64'h676e6172_2d656761,
        64'h746c6f76_0079636e,
        64'h65757165_72662d78,
        64'h616d2d69_7073006f,
        64'h69746172_2d6b6373,
        64'h2c786e6c_78007374,
        64'h69622d72_6566736e,
        64'h6172742d_6d756e2c,
        64'h786e6c78_00737469,
        64'h622d7373_2d6d756e,
        64'h2c786e6c_78007473,
        64'h6978652d_6f666966,
        64'h2c786e6c_7800796c,
        64'h696d6166_2c786e6c,
        64'h78006874_6469772d,
        64'h6f692d67_65720074,
        64'h66696873_2d676572,
        64'h00737470_75727265,
        64'h746e6900_746e6572,
        64'h61702d74_70757272,
        64'h65746e69_00646565,
        64'h70732d74_6e657272,
        64'h75630076_65646e2c,
        64'h76637369_72007974,
        64'h69726f69_72702d78,
        64'h616d2c76_63736972,
        64'h0073656d_616e2d67,
        64'h65720064_65646e65,
        64'h7478652d_73747075,
        64'h72726574_6e690073,
        64'h65676e61_7200656c,
        64'h646e6168_702c7875,
        64'h6e696c00_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h00687461_702d7475,
        64'h6f647473_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h02000000_02000000,
        64'h03000000_bb000000,
        64'h04000000_03000000,
        64'h03000000_b5000000,
        64'h04000000_03000000,
        64'h01000000_67000000,
        64'h04000000_03000000,
        64'h00000000_7968702d,
        64'h74656e72_65687465,
        64'h5b000000_0d000000,
        64'h03000000_00000000,
        64'h35313963_2e633130,
        64'h3064692d_7968702d,
        64'h74656e72_65687465,
        64'h1b000000_19000000,
        64'h03000000_00003040,
        64'h7968702d_74656e72,
        64'h65687465_01000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_6f69646d,
        64'h01000000_00000000,
        64'h64692d69_696d6772,
        64'ha2020000_09000000,
        64'h03000000_01000000,
        64'h94020000_04000000,
        64'h03000000_00000000,
        64'h82020000_04000000,
        64'h03000000_01000000,
        64'h70020000_04000000,
        64'h03000000_04000000,
        64'h5c020000_04000000,
        64'h03000000_01000000,
        64'h4a020000_04000000,
        64'h03000000_00657469,
        64'h6c74656e_72656874,
        64'h655f6978_615f786e,
        64'h6c785f69_3c020000,
        64'h18000000_03000000,
        64'h01000000_2a020000,
        64'h04000000_03000000,
        64'h00000000_0b020000,
        64'h04000000_03000000,
        64'h01000000_ef010000,
        64'h04000000_03000000,
        64'h01000000_e3010000,
        64'h04000000_03000000,
        64'h00000100_00000000,
        64'h00000030_00000000,
        64'h67000000_10000000,
        64'h03000000_03000000,
        64'hd8010000_04000000,
        64'h03000000_00002201,
        64'h00350a00_c6010000,
        64'h06000000_03000000,
        64'h00000000_03000000,
        64'h25010000_08000000,
        64'h03000000_02000000,
        64'h14010000_04000000,
        64'h03000000_006b726f,
        64'h7774656e_5b000000,
        64'h08000000_03000000,
        64'h0000612e_30302e31,
        64'h2d657469_6c74656e,
        64'h72656874_652d7370,
        64'h782c786e_6c780030,
        64'h2e332d65_74696c74,
        64'h656e7265_6874652d,
        64'h6978612c_786e6c78,
        64'h1b000000_37000000,
        64'h03000000_00000030,
        64'h30303030_30303340,
        64'h74656e72_65687465,
        64'h01000000_02000000,
        64'h02000000_bb010000,
        64'h00000000_03000000,
        64'he40c0000_e40c0000,
        64'hac010000_08000000,
        64'h03000000_20bcbe00,
        64'h9a010000_04000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00000000,
        64'h746f6c73_2d697073,
        64'h2d636d6d_1b000000,
        64'h0d000000_03000000,
        64'h00000030_40636d6d,
        64'h01000000_04000000,
        64'h8b010000_04000000,
        64'h03000000_08000000,
        64'h74010000_04000000,
        64'h03000000_01000000,
        64'h63010000_04000000,
        64'h03000000_01000000,
        64'h53010000_04000000,
        64'h03000000_00377865,
        64'h746e696b_47010000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h00000020_00000000,
        64'h67000000_10000000,
        64'h03000000_02000000,
        64'h02000000_25010000,
        64'h08000000_03000000,
        64'h02000000_14010000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00612e30_302e322d,
        64'h6970732d_7370782c,
        64'h786e6c78_00622e30,
        64'h302e322d_6970732d,
        64'h7370782c_786e6c78,
        64'h1b000000_28000000,
        64'h03000000_00000000,
        64'h30303030_30303032,
        64'h40697073_2d737078,
        64'h01000000_02000000,
        64'h04000000_3a010000,
        64'h04000000_03000000,
        64'h02000000_30010000,
        64'h04000000_03000000,
        64'h01000000_25010000,
        64'h04000000_03000000,
        64'h02000000_14010000,
        64'h04000000_03000000,
        64'h00c20100_06010000,
        64'h04000000_03000000,
        64'h80f0fa02_4b000000,
        64'h04000000_03000000,
        64'h00100000_00000000,
        64'h00000010_00000000,
        64'h67000000_10000000,
        64'h03000000_00303537,
        64'h3631736e_1b000000,
        64'h08000000_03000000,
        64'h00000030_30303030,
        64'h30303140_74726175,
        64'h01000000_02000000,
        64'h006c6f72_746e6f63,
        64'hde000000_08000000,
        64'h03000000_00100000,
        64'h00000000_00000000,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'hffff0000_01000000,
        64'hca000000_08000000,
        64'h03000000_00333130,
        64'h2d677562_65642c76,
        64'h63736972_1b000000,
        64'h10000000_03000000,
        64'h00003040_72656c6c,
        64'h6f72746e_6f632d67,
        64'h75626564_01000000,
        64'h02000000_02000000,
        64'hbb000000_04000000,
        64'h03000000_02000000,
        64'hb5000000_04000000,
        64'h03000000_03000000,
        64'hfb000000_04000000,
        64'h03000000_07000000,
        64'he8000000_04000000,
        64'h03000000_00000004,
        64'h00000000_0000000c,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h09000000_01000000,
        64'h0b000000_01000000,
        64'hca000000_10000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h00306369_6c702c76,
        64'h63736972_1b000000,
        64'h0c000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_00000000,
        64'h04000000_03000000,
        64'h00000000_30303030,
        64'h30306340_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_02000000,
        64'h006c6f72_746e6f63,
        64'hde000000_08000000,
        64'h03000000_00000c00,
        64'h00000000_00000002,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h07000000_01000000,
        64'h03000000_01000000,
        64'hca000000_10000000,
        64'h03000000_00000000,
        64'h30746e69_6c632c76,
        64'h63736972_1b000000,
        64'h0d000000_03000000,
        64'h00000030_30303030,
        64'h30324074_6e696c63,
        64'h01000000_c3000000,
        64'h00000000_03000000,
        64'h00007375_622d656c,
        64'h706d6973_00636f73,
        64'h2d657261_622d656e,
        64'h61697261_2c687465,
        64'h1b000000_1f000000,
        64'h03000000_02000000,
        64'h0f000000_04000000,
        64'h03000000_02000000,
        64'h00000000_04000000,
        64'h03000000_00636f73,
        64'h01000000_02000000,
        64'h00000008_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h01000000_bb000000,
        64'h04000000_03000000,
        64'h01000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00007573_63616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'h40787d01_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30314074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h10090000_ab020000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h48090000_38000000,
        64'hf30b0000_edfe0dd0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'ha0018402_17c58593,
        64'h00000597_01f41413,
        64'h0010041b_e911d13f,
        64'hf0ef057e_65a14505,
        64'hef6ff0ef_d9450513,
        64'h00001517_ed0ff0ef,
        64'he4061141_b38df0cf,
        64'hf0ef07a5_05130000,
        64'h1517bbd9_df450513,
        64'h00001517_fa4ff0ef,
        64'h8526f28f_f0efed65,
        64'h05130000_1517f34f,
        64'hf0efeca5_05130000,
        64'h1517bbfd_e1c50513,
        64'h00001517_fccff0ef,
        64'h8526f50f_f0efefe5,
        64'h05130000_1517f5cf,
        64'hf0efef25_05130000,
        64'h1517c929_84aac69f,
        64'hf0ef8556_865e020b,
        64'h2583f78f_f0ef0ce5,
        64'h05130000_1517f384,
        64'h9de30809_0913080a,
        64'h0993f90f_f0ef2485,
        64'he7050513_00001517,
        64'hff3a1be3_867ff0ef,
        64'h0a05000a_4503facf,
        64'hf0ef0f25_05130000,
        64'h151783bf_f0ef0109,
        64'h3503fc0f_f0ef0f65,
        64'h05130000_151784ff,
        64'hf0ef0089_3503fd4f,
        64'hf0ef0fa5_05130000,
        64'h1517863f_f0effb89,
        64'h8a130009_3503fecf,
        64'hf0ef1025_05130000,
        64'h1517ff2a_1be38c1f,
        64'hf0ef0a05_000a4503,
        64'hf9098a13_80bff0ef,
        64'h10050513_00001517,
        64'hff9a19e3_8dfff0ef,
        64'h0a050007_c503014d,
        64'h07b34a01_82bff0ef,
        64'hf8098d13_10450513,
        64'h00001517_8ffff0ef,
        64'h0ff4f513_843ff0ef,
        64'h10050513_00001517,
        64'h4c114cc1_10051b63,
        64'h02010913_08010993,
        64'h84aa8b0a_d5fff0ef,
        64'h850a4605_71010489,
        64'h2583871f_f0eff4e5,
        64'h05130000_15178bff,
        64'hf0ef4556_883ff0ef,
        64'h12050513_00001517,
        64'h8d1ff0ef_4546895f,
        64'hf0ef1125_05130000,
        64'h1517923f_f0ef6526,
        64'h8a7ff0ef_10450513,
        64'h00001517_935ff0ef,
        64'h75028b9f_f0ef1065,
        64'h05130000_1517947f,
        64'hf0ef6562_8cbff0ef,
        64'h10050513_00001517,
        64'h919ff0ef_45528ddf,
        64'hf0ef1025_05130000,
        64'h151792bf_f0ef4542,
        64'h8efff0ef_10450513,
        64'h00001517_93dff0ef,
        64'h4532901f_f0ef1065,
        64'h05130000_151794ff,
        64'hf0ef4522_913ff0ef,
        64'h10850513_00001517,
        64'h9a1ff0ef_6502925f,
        64'hf0ef10a5_05130000,
        64'h1517931f_f0ef0f65,
        64'h05130000_1517bf51,
        64'h54f9941f_f0ef01e5,
        64'h05130000_15179cff,
        64'hf0ef8526_953ff0ef,
        64'h10050513_00001517,
        64'h95fff0ef_0f450513,
        64'h00001517_c90584aa,
        64'h890ae6df_f0ef850a,
        64'h45854605_710197df,
        64'hf0ef0fa5_05130000,
        64'h15178082_61256d02,
        64'h6ca26c42_6be27b02,
        64'h7aa27a42_79e26906,
        64'h64a66446_852660e6,
        64'hfa040113_54fd9adf,
        64'hf0ef1025_05130000,
        64'h1517c90d_e1bff0ef,
        64'h8bae8aaa_1080e06a,
        64'he466e862_f05af852,
        64'hfc4ee0ca_e4a6ec86,
        64'hec5ef456_e8a2711d,
        64'hbfe15479_80826169,
        64'h6baa6b4a_6aea7a0a,
        64'h79aa794a_74ea640e,
        64'h60ae8522_c7bff0ef,
        64'hc87ff0ef_45314581,
        64'h46054401_f89046e3,
        64'h20090913_14fda15f,
        64'hf0ef1625_05130000,
        64'h1517e799_0364e7b3,
        64'h04899463_90412981,
        64'h14428c49_cb3ff0ef,
        64'h90410305_14130085,
        64'h151bcc1f_f0effd24,
        64'h1ae30404_0413ff7a,
        64'h17e389aa_f11ff0ef,
        64'h0a05854e_0007c583,
        64'h014407b3_04000b93,
        64'h4a01c65f_f0ef850a,
        64'h04000593_86224981,
        64'hff551ee3_cfbff0ef,
        64'he0090413_3e800b13,
        64'h0fe00a93_20090913,
        64'h90811482_bff5d15f,
        64'hf0efc501_d23ff0ef,
        64'h454985a2_0ff67613,
        64'h00166613_0015161b,
        64'hf53ff0ef_0ff47593,
        64'hf5bff0ef_0ff5f593,
        64'h0084559b_f67ff0ef,
        64'h0ff5f593_0104559b,
        64'hf73ff0ef_45010184,
        64'h559bfee7_9be30785,
        64'h00c68023_00f106b3,
        64'h08000713_567d4781,
        64'h842e892a_e55ee95a,
        64'hed56f152_f54ee586,
        64'h84b2f94a_fd26e1a2,
        64'h71558082_91411542,
        64'h8d3d8ff9_0057979b,
        64'h17016709_0107d79b,
        64'h0105179b_4105551b,
        64'h0105151b_8d2d00c5,
        64'h95138da9_893d0045,
        64'hd51b8da9_91411542,
        64'h8d5d0522_0085579b,
        64'h808207f5_75138d2d,
        64'h00451593_8d2d8d3d,
        64'h0045d51b_0075d79b,
        64'h8de98082_0141853e,
        64'h640260a2_57f5e111,
        64'h4781f89f_f0efc511,
        64'h57f9efbf_f0efc911,
        64'h57fdeb7f_f0effc6d,
        64'he07ff0ef_347d4429,
        64'hb8fff0ef_2c450513,
        64'h00001517_c89ff0ef,
        64'he022e406_11418082,
        64'h61050015_351364a2,
        64'h644260e2_0004051b,
        64'hfc940ce3_e3bff0ef,
        64'heb3ff0ef_2ec50513,
        64'h00001517_85aa842a,
        64'he57ff0ef_02900513,
        64'h400005b7_07700613,
        64'hfbdff0ef_4485e822,
        64'hec06e426_11018082,
        64'h01410015_3513157d,
        64'h640260a2_0004051b,
        64'hef3ff0ef_32650513,
        64'h85a20000_1517e8df,
        64'hf0ef842a_e9bff0ef,
        64'he022e406_03700513,
        64'h45810650_06131141,
        64'h80826105_690264a2,
        64'h644260e2_00153513,
        64'hf5650513_0004051b,
        64'h01249863_88bd00f9,
        64'h1b634501_4785ecdf,
        64'hf0efed1f_f0ef842a,
        64'hed7ff0ef_84aaeddf,
        64'hf0efee1f_f0efee5f,
        64'hf0ef892a_ef3ff0ef,
        64'he04ae426_e822ec06,
        64'h45211aa0_05930870,
        64'h06131101_bfcd4501,
        64'h80826105_690264a2,
        64'h644260e2_4505f89f,
        64'hf0ef4585_3b450513,
        64'h00001517_fe9915e3,
        64'hc00df29f_f0ef892a,
        64'h347df39f_f0ef4501,
        64'h45810950_06134485,
        64'h71040413_e04aec06,
        64'he4266409_e8221101,
        64'hccfff06f_61053ae5,
        64'h05130000_151760e2,
        64'h6442da5f_f0ef852e,
        64'h65a2ce9f_f0ef3f65,
        64'h05130000_1517cf5f,
        64'hf0ef8522_cfbff0ef,
        64'he42eec06_3fc50513,
        64'h00001517_842ae822,
        64'h11018082_614564e2,
        64'h740270a2_f47d147d,
        64'h0007d463_4187d79b,
        64'h0185179b_fabff0ef,
        64'heb5ff0ef_85320640,
        64'h04136622_ec1ff0ef,
        64'h0ff47513_ec9ff0ef,
        64'h0ff57513_0084551b,
        64'hed5ff0ef_0ff57513,
        64'h0104551b_ee1ff0ef,
        64'h0184551b_ee9ff0ef,
        64'h0404e513_febff0ef,
        64'h84aa842e_ec26f022,
        64'he432f406_7179f03f,
        64'hf06f0ff0_05138082,
        64'h557db7d9_00d70023,
        64'h078500f6_073306c8,
        64'h2683ff69_8b055178,
        64'hb77dd6b8_07850007,
        64'h470300f5_07338082,
        64'h4501d3b8_4719dbb8,
        64'h577d2000_07b702b6,
        64'he1630007_869b2000,
        64'h08372000_0537fff5,
        64'h8b85537c_20000737,
        64'hd3b82000_07b71060,
        64'h0713fff5_37fd0001,
        64'h03200793_04b76163,
        64'h0007871b_47812000,
        64'h06b7dbb8_57792000,
        64'h07b706b7_ee631000,
        64'h07938082_610564a2,
        64'hd3b84719_dbb86442,
        64'h60e20ff4_7513577d,
        64'h200007b7_e23ff0ef,
        64'h50050513_00001517,
        64'heb1ff0ef_91011502,
        64'h4088e39f_f0ef51e5,
        64'h05130000_1517e395,
        64'h8b852401_53fc57e0,
        64'hff658b05_06478493,
        64'h53f8d3b8_10600713,
        64'h200007b7_fff537fd,
        64'h00010640_0793d7a8,
        64'hdbb85779_e426e822,
        64'hec062000_07b71101,
        64'he7fff06f_610554e5,
        64'h05130000_151764a2,
        64'h60e26442_d03c4799,
        64'he97ff0ef_57450513,
        64'h00001517_f25ff0ef,
        64'h91010204_95132481,
        64'heafff0ef_56c50513,
        64'h00001517_5064d03c,
        64'h16600793_ec3ff0ef,
        64'h5a050513_00001517,
        64'hf51ff0ef_91010204,
        64'h95132481_edbff0ef,
        64'h59850513_00001517,
        64'h5064d03c_10400793,
        64'h20000437_fff537fd,
        64'h000147a9_c3b84729,
        64'h200007b7_f03ff0ef,
        64'he426e822_ec065b85,
        64'h05131101_00001517,
        64'h80822501_41088082,
        64'hc10c8082_610560e2,
        64'hee1ff0ef_00914503,
        64'hee9ff0ef_00814503,
        64'hf55ff0ef_ec06002c,
        64'h11018082_61456942,
        64'h64e27402_70a2fe94,
        64'h10e3f0bf_f0ef0091,
        64'h4503f13f_f0ef3461,
        64'h00814503_f81ff0ef,
        64'h0ff57513_002c0089,
        64'h553354e1_03800413,
        64'h892af406_e84aec26,
        64'hf0227179_80826145,
        64'h694264e2_740270a2,
        64'hfe9410e3_f4dff0ef,
        64'h00914503_f55ff0ef,
        64'h34610081_4503fc3f,
        64'hf0ef0ff5_7513002c,
        64'h0089553b_54e14461,
        64'h892af406_e84aec26,
        64'hf0227179_808200f5,
        64'h80230007_c78300e5,
        64'h80a397aa_81110007,
        64'h4703973e_00f57713,
        64'h98078793_00001797,
        64'hb7f50405_fa5ff0ef,
        64'h80820141_640260a2,
        64'he5090004_4503842a,
        64'he406e022_11418082,
        64'h00e78823_02000713,
        64'h00e78423_fc700713,
        64'h00e78623_470d0007,
        64'h822300e7_8023476d,
        64'h00e78623_f8000713,
        64'h00078223_100007b7,
        64'h808200a7_0023dfe5,
        64'h0207f793_01474783,
        64'h10000737_80820205,
        64'h75130147_c5031000,
        64'h07b78082_00054503,
        64'h808200b5_00238082,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00048067_01f49493,
        64'h0010049b_b8458593,
        64'h00001597_f1402573,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'hfe091ee3_0004a903,
        64'h00092023_00990933,
        64'h00291913_f1402973,
        64'h020004b7_fe090ae3,
        64'h00897913_34402973,
        64'h10500073_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_0124a023,
        64'h00100913_020004b7,
        64'h241000ef_01a11113,
        64'h0210011b_03249663,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
